constant_inst : constant PORT MAP (
		result	 => result_sig
	);
