const1_inst : const1 PORT MAP (
		result	 => result_sig
	);
